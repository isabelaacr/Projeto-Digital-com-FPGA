-- Faça um circuito que tenha 5 bits de entrada e 3 saídas.
-- A lógica do circuito é dada por uma tabela verdade única (gerada por você e diferente de todos os demais colegas de aula).
-- Faça a programação, que implemente o circuito projetado, e faça também o test bench para fazer a simulação do circuito, explorando no mínimo 15 das 32 possibilidades da entrada.
-- Faça um relatório para apresentação do projeto, bem como a simulação do mesmo.

