library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity principal is
    Port (
        numero : in integer range 0 to 9;
        d      : out STD_LOGIC_VECTOR(6 downto 0);
        sel    : out STD_LOGIC_VECTOR(3 downto 0)
    );
end principal;

architecture Behavioral of principal is

    component disp
        Port (
            n : in integer range 0 to 9;
            d : out STD_LOGIC_VECTOR(6 downto 0)
        );
    end component;

begin

    sel <= "1110";

    ul: disp port map (
        n => numero,
        d => d
    );

end Behavioral;
